`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/18/2016 03:02:01 PM
// Design Name: 
// Module Name: char_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module char_rom(
   output [15:0] DO,     // Output data, width defined by READ_WIDTH parameter
   input [10:0] ADDR,   // Input address, width defined by read/write port depth
   input CLK,           // 1-bit input clock
   input [15:0] DI,      // Input data port, width defined by WRITE_WIDTH parameter
   input EN,            // 1-bit input RAM enable
   input REGCE,         // 1-bit input output register enable
   input RST,           // 1-bit input reset
   input [1:0] WE             // Input write enable, width defined by write port depth
   );
    
// BRAM_SINGLE_MACRO: Single Port RAM
//                    Artix-7
// Xilinx HDL Language Template, version 2016.2

/////////////////////////////////////////////////////////////////////
//  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            //
// WRITE_WIDTH |           | WRITE Depth |            |  WE Width  //
// ============|===========|=============|============|============//
//    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   //
//    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   //
//    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   //
//    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   //
//    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   //
//     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   //
//     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   //
//     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   //
//     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   //
//       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   //
//       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   //
//       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   //
//       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   //
/////////////////////////////////////////////////////////////////////

BRAM_SINGLE_MACRO #(
   .BRAM_SIZE("36Kb"), // Target BRAM, "18Kb" or "36Kb" 
   .DEVICE("7SERIES"), // Target Device: "7SERIES" 
   .DO_REG(0), // Optional output register (0 or 1)
   .INIT(9'h000000000), // Initial values on output port
   .INIT_FILE ("NONE"),
   .WRITE_WIDTH(16), // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
   .READ_WIDTH(16),  // Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
   .SRVAL(9'h0), // Set/Reset value for port output
   .WRITE_MODE("WRITE_FIRST"), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE" 
   .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INIT_21(256'h0000000003000300030003000300030003000300030000000300030000000000),
   .INIT_22(256'h0000000006600660066006600000000000000000000000000000000000000000),
   .INIT_23(256'h000000000360036006C03FF03FF006C00D803FF03FF00D801B001B0000000000),
   .INIT_24(256'h00000100038007C00D600D000F00078003C001E00D600D6007C0038001000000),
   .INIT_25(256'h000000003C1866306630666066C03CC0019E01B30333033306330C1E00000000),
   .INIT_26(256'h0000000007C00FE00C600C6007C007800D9019D818F018780FFC078800000000),
   .INIT_27(256'h0000000001800180018001800000000000000000000000000000000000000000),
   .INIT_28(256'h0000018003000300060006000600060006000600060003000300018000000000),
   .INIT_29(256'h0000060003000300018001800180018001800180018003000300060000000000),
   .INIT_2A(256'h00000000000000000380038033983FF807C007C00EE01C700440000000000000),
   .INIT_2B(256'h0000000000000000000000C000C000C007F807F800C000C000C0000000000000),
   .INIT_2C(256'h0000000000000000000000000000000000000000030003000100010002000000),
   .INIT_2D(256'h0000000000000000000000000000000003E003E0000000000000000000000000),
   .INIT_2E(256'h0000000000000000000000000000000000000000000003000300000000000000),
   .INIT_2F(256'h000000000060006000C000C000C000C001800180018001800300030000000000),
   .INIT_30(256'h0000000003C007E00E700C300C300C300C300C300C300E7007E003C000000000),
   .INIT_31(256'h000000000180038007800D800980018001800180018001800180018000000000),
   .INIT_32(256'h0000000003C007E00E300C300030006000E001C0038006000FF00FF000000000),
   .INIT_33(256'h0000000003E007F00E30003001E001E0007000300C300E7007E003C000000000),
   .INIT_34(256'h00000000006000E000E001E00360036006600C600FF00FF00060006000000000),
   .INIT_35(256'h0000000007E007E006000C000FC00FE00C7000300C300E7007E003C000000000),
   .INIT_36(256'h0000000003E007F006300C000DC00FE00E700C300C30063007E003C000000000),
   .INIT_37(256'h000000000FF00FF0006000C000C0018001800180038003000300030000000000),
   .INIT_38(256'h0000000003C007E00C300C300C3007E007E00C300C300C3007E003C000000000),
   .INIT_39(256'h0000000003C007E00C600C300C300E7007F003B000300C600FE007C000000000),
   .INIT_3A(256'h0000000000000180018000000000000000000000018001800000000000000000),
   .INIT_3B(256'h0000000000000180018000000000000000000000018001800080008001000000),
   .INIT_3C(256'h0000000000000000002000E003C00F001C000F0003C000E00020000000000000),
   .INIT_3D(256'h00000000000000001FF01FF0000000001FF01FF0000000000000000000000000),
   .INIT_3E(256'h000000000000000008000E00078001E0007001E007800E000800000000000000),
   .INIT_3F(256'h0000000003C007E00E300C30007000E001C00180018000000180018000000000),
   .INIT_40(256'h000007C00C30137817E82CC82CC82CC82FD026E01008081007E0000000000000),
   .INIT_41(256'h000000000380038006C006C006C00C600C600FE01FF018301830301800000000),
   .INIT_42(256'h000000001FE01FF01830183018301FE01FF01818181818181FF01FE000000000),
   .INIT_43(256'h0000000003E00FF00C381C1018001800180018001C100C380FF003E000000000),
   .INIT_44(256'h000000001FC01FF0183018181818181818181818181818301FF01FC000000000),
   .INIT_45(256'h000000000FF80FF80C000C000C000FF80FF80C000C000C000FF80FF800000000),
   .INIT_46(256'h000000000FF00FF00C000C000C000FE00FE00C000C000C000C000C0000000000),
   .INIT_47(256'h0000000007E01FF0183838103000300030F830F8381818381FF807E000000000),
   .INIT_48(256'h00000000181818181818181818181FF81FF81818181818181818181800000000),
   .INIT_49(256'h0000000001800180018001800180018001800180018001800180018000000000),
   .INIT_4A(256'h00000000003000300030003000300030003000300C300E7007E003C000000000),
   .INIT_4B(256'h0000000018181830186018C019801BC01EC01C60187018301818181800000000),
   .INIT_4C(256'h000000000C000C000C000C000C000C000C000C000C000C000FF00FF000000000),
   .INIT_4D(256'h00000000383838383C783C78345836D836D836D8339833983398311800000000),
   .INIT_4E(256'h0000000018181C181E181E181B181998199818D8187818781838181800000000),
   .INIT_4F(256'h0000000007C01FF0183030183018301830183018301818301FF007C000000000),
   .INIT_50(256'h000000000FE00FF00C380C180C380FF00FE00C000C000C000C000C0000000000),
   .INIT_51(256'h0000000007C01FF018303018301830183018301831B818F01FF007B000180000),
   .INIT_52(256'h000000001FE01FF01838181818381FF01FC018E0187018301838181C00000000),
   .INIT_53(256'h0000000003E007F00E380C180F0007E001F000380C180E3807F003E000000000),
   .INIT_54(256'h000000001FF81FF8018001800180018001800180018001800180018000000000),
   .INIT_55(256'h000000001818181818181818181818181818181818181C380FF007E000000000),
   .INIT_56(256'h0000000030181830183018300C600C600EE006C006C003800380038000000000),
   .INIT_57(256'h0000000031C631C631C61B6C1B6C1B6C1B6C1B6C0E380E380E380E3800000000),
   .INIT_58(256'h0000000018301C700C6006C007C00380038007C006C00C601C70183000000000),
   .INIT_59(256'h0000000018181C380C300660066003C001800180018001800180018000000000),
   .INIT_5A(256'h0000000007F807F80030006000E000C001800380030006000FF80FF800000000),
   .INIT_5B(256'h000003C003C0030003000300030003000300030003000300030003C003C00000),
   .INIT_5C(256'h0000000003000300018001800180018000C000C000C000C00060006000000000),
   .INIT_5D(256'h000003C003C000C000C000C000C000C000C000C000C000C000C003C003C00000),
   .INIT_5E(256'h0000018003C003C00660066006600C3000000000000000000000000000000000),
   .INIT_5F(256'h0000000000000000000000000000000000000000000000000000FFFFFFFF0000),
   .INIT_60(256'h00000000018000C0000000000000000000000000000000000000000000000000),
   .INIT_61(256'h000000000000000007C00FE00C6001E007E00E600C600FE007B0000000000000),
   .INIT_62(256'h00000C000C000C000DC00FE00E700C300C300C300E700FE00DC0000000000000),
   .INIT_63(256'h000000000000000003C007E00E600C000C000C000E6007E003C0000000000000),
   .INIT_64(256'h000000300030003003B007F00E700C300C300C300E7007F003B0000000000000),
   .INIT_65(256'h0000000000000000038007C00C600FE00FE00C000E6007C00380000000000000),
   .INIT_66(256'h000003C007C006000F800F800600060006000600060006000600000000000000),
   .INIT_67(256'h00000000000007600FE01CE01860186018601CE00FE0076018601FE00FC00000),
   .INIT_68(256'h00000C000C000C000DE00FF00E300C300C300C300C300C300C30000000000000),
   .INIT_69(256'h0000000001800180000001800180018001800180018001800180000000000000),
   .INIT_6A(256'h0000000001800180000001800180018001800180018001800180018007800700),
   .INIT_6B(256'h00000C000C000C000C600CC00D800F800FC00EC00CC00C600C60000000000000),
   .INIT_6C(256'h0000018001800180018001800180018001800180018001800180000000000000),
   .INIT_6D(256'h000000000000000037383FFC39CC318C318C318C318C318C318C000000000000),
   .INIT_6E(256'h00000000000000000DE00FF00E300C300C300C300C300C300C30000000000000),
   .INIT_6F(256'h000000000000000003C007E00E700C300C300C300E7007E003C0000000000000),
   .INIT_70(256'h00000000000000000DC00FE00E700C300C300C300E700FE00DC00C000C000C00),
   .INIT_71(256'h000000000000000003B007F00E700C300C300C300E7007F003B0003000300030),
   .INIT_72(256'h0000000000000000037003F00380030003000300030003000300000000000000),
   .INIT_73(256'h000000000000000007C00FE00C600F0007C000E00C600FE007C0000000000000),
   .INIT_74(256'h000001000300030007C007C00300030003000300030003C001C0000000000000),
   .INIT_75(256'h00000000000000000C300C300C300C300C300C300C700FF007B0000000000000),
   .INIT_76(256'h000000000000000006300630063003600360036001C001C001C0000000000000),
   .INIT_77(256'h000000000000000031C631C619CC1B6C1B6C1B6C0E380E380E38000000000000),
   .INIT_78(256'h000000000000000006300770036001C001C001C0036007700630000000000000),
   .INIT_79(256'h00000000000000000C180C18063006300360036003E001C001C0018007800700),
   .INIT_7A(256'h000000000000000003F803F80030007000E001C0018003F803F8000000000000),
   .INIT_7B(256'h01C003C003000300030003000E000E000300030003000300030003C001C00000),
   .INIT_7C(256'h0180018001800180018001800180018001800180018001800180018001800180),
   .INIT_7D(256'h038003C000C000C000C000C00070007000C000C000C000C000C003C003800000),
   .INIT_7E(256'h0000000007880FF808F000000000000000000000000000000000000000000000),
   .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
   
   // The next set of INITP_xx are for the parity bits
   .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
   
   // The next set of INIT_xx are valid when configured as 36Kb
   .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
   .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)
) BRAM_SINGLE_MACRO_inst (
   .DO(DO),       // Output data, width defined by READ_WIDTH parameter
   .ADDR(ADDR),   // Input address, width defined by read/write port depth
   .CLK(CLK),     // 1-bit input clock
   .DI(DI),       // Input data port, width defined by WRITE_WIDTH parameter
   .EN(EN),       // 1-bit input RAM enable
   .REGCE(REGCE), // 1-bit input output register enable
   .RST(RST),     // 1-bit input reset
   .WE(WE)        // Input write enable, width defined by write port depth
);

// End of BRAM_SINGLE_MACRO_inst instantiation
                

endmodule


